`include "./../conf/conf.v"

module register_file(
    input [4:0] rx,

    output [ISA_WIDTH-1:0] word_o
);



endmodule
